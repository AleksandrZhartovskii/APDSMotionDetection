library ieee;
use ieee.std_logic_1164.all;

entity frequency_controller is

    port (
        clk_in  : in  std_logic;
        clk_out : out std_logic
    );

end frequency_controller;

architecture rtl of frequency_controller is     
begin



end rtl;
